library verilog;
use verilog.vl_types.all;
entity FF_DUT is
end FF_DUT;
