library verilog;
use verilog.vl_types.all;
entity Counter_DUT is
end Counter_DUT;
