// ---------------------------   T Flip Flop   ------------------------------- //
module FF ( clk , reset , D , Q ) ;
// -------------------------- Inputs Declarations ---------------------------- //
input clk , D, reset ;
// ------------------------- Outputs Declarations ---------------------------- //
output Q ;
// ---------------------------- Reg Declarations ----------------------------- //
reg Q ;
always @( posedge clk or posedge reset)
begin
  if(reset)
	  Q <= 0 ;
  else
	  Q <= ~D ;
end

endmodule
// ----------------------------- End of File --------------------------------- //
// --------------------------------------------------------------------------- //
