library verilog;
use verilog.vl_types.all;
entity sevenSegments_DUT is
end sevenSegments_DUT;
