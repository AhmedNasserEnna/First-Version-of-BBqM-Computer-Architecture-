library verilog;
use verilog.vl_types.all;
entity Display_DUT is
end Display_DUT;
