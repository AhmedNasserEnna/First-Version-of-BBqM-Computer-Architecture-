library verilog;
use verilog.vl_types.all;
entity ROM_DUT is
end ROM_DUT;
