library verilog;
use verilog.vl_types.all;
entity BBqM_DUT is
end BBqM_DUT;
