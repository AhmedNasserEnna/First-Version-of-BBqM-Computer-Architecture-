library verilog;
use verilog.vl_types.all;
entity clock_divider_DUT is
end clock_divider_DUT;
