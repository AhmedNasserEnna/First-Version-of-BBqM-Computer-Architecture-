library verilog;
use verilog.vl_types.all;
entity UpDown_Counter_FSM_DUT is
end UpDown_Counter_FSM_DUT;
